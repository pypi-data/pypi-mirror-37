dimensions:
	dim0 = 1 ;
	lat = 2 ;
	lon = 2 ;
variables:
	double temp(lon, lat) ;
		temp:standard_name = "surface_temperature" ;
		temp:units = "K" ;
	int64 lon(lon) ;
		lon:axis = "X" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
	int64 lat(lat) ;
		lat:units = "degree_north" ;
	double temp2(dim0, lon, lat) ;
		temp2:long_name = "Something Random" ;
		temp2:units = "K" ;
	int64 dim0(dim0) ;
		dim0:long_name = "Rnd Coordinate" ;

// global attributes:
		:Conventions = "CF-1.5" ;
}
